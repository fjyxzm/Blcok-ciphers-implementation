`timescale 1ns/1ns
`define    N      63

module MixColumn(c,b);   //c=a*b
    input  [`N:0] b;
    output [`N:0] c;
    
    reg    [`N:0] a;
    wire   [`N:0] c;
    
    initial  begin
	  a[63:60]=4; a[59:56]= 1; a[55:52]= 2; a[51:48]= 2;
	  a[47:44]=8; a[43:40]= 6; a[39:36]= 5; a[35:32]= 6;
	  a[31:28]=11;a[27:24]=14; a[23:20]=10; a[19:16]= 9;
	  a[15:12]= 2;a[11: 8]= 2; a[ 7: 4]=15; a[ 3: 0]=11;
    end  
    
    
    FieldMutilSum sum00(c[63:60],a[63:60],a[59:56],a[55:52],a[51:48],
                                b[63:60],b[47:44],b[31:28],b[15:12]);
    FieldMutilSum sum01(c[59:56],a[63:60],a[59:56],a[55:52],a[51:48],
                                b[59:56],b[43:40],b[27:24],b[11:8]);
    FieldMutilSum sum02(c[55:52],a[63:60],a[59:56],a[55:52],a[51:48],
                                b[55:52],b[39:36],b[23:20],b[7:4]);
    FieldMutilSum sum03(c[51:48],a[63:60],a[59:56],a[55:52],a[51:48],
                                b[51:48],b[35:32],b[19:16],b[3:0]);
                         
    FieldMutilSum sum10(c[47:44],a[47:44],a[43:40],a[39:36],a[35:32],
                                b[63:60],b[47:44],b[31:28],b[15:12]);
    FieldMutilSum sum11(c[43:40],a[47:44],a[43:40],a[39:36],a[35:32],
                                b[59:56],b[43:40],b[27:24],b[11:8]);
    FieldMutilSum sum12(c[39:36],a[47:44],a[43:40],a[39:36],a[35:32],
                                b[55:52],b[39:36],b[23:20],b[7:4]);
    FieldMutilSum sum13(c[35:32],a[47:44],a[43:40],a[39:36],a[35:32],
                                b[51:48],b[35:32],b[19:16],b[3:0]);
                         
    FieldMutilSum sum20(c[31:28],a[31:28],a[27:24],a[23:20],a[19:16],
                                b[63:60],b[47:44],b[31:28],b[15:12]);
    FieldMutilSum sum21(c[27:24],a[31:28],a[27:24],a[23:20],a[19:16],
                                b[59:56],b[43:40],b[27:24],b[11:8]);
    FieldMutilSum sum22(c[23:20],a[31:28],a[27:24],a[23:20],a[19:16],
                                b[55:52],b[39:36],b[23:20],b[7:4]);
    FieldMutilSum sum23(c[19:16],a[31:28],a[27:24],a[23:20],a[19:16],
                                b[51:48],b[35:32],b[19:16],b[3:0]);
                         
    
    FieldMutilSum sum30(c[15:12],a[15:12],a[11:8],a[7:4],a[3:0],
                                b[63:60],b[47:44],b[31:28],b[15:12]);
    FieldMutilSum sum31(c[11:8], a[15:12],a[11:8],a[7:4],a[3:0],
                                b[59:56],b[43:40],b[27:24],b[11:8]);
    FieldMutilSum sum32(c[7:4],  a[15:12],a[11:8],a[7:4],a[3:0],
                                b[55:52],b[39:36],b[23:20],b[7:4]);
    FieldMutilSum sum33(c[3:0],  a[15:12],a[11:8],a[7:4],a[3:0],
                                b[51:48],b[35:32],b[19:16],b[3:0]);
    
 endmodule 